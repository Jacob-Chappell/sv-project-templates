`timescale 1ns / 10ps

// Created for ${For} in the ${PROJECT_NAME}
// Description: ${Description}

module ${NAME} #(
    
) (
    #if(${Is_Clocked}==true)input clk, n_rst, // Clock period = ${Clock_Period}#end
);

    

endmodule
