`timescale 1ns / 10ps

// Created for ${ORGANIZATION} in the ${PROJECT_NAME} project

module ${MOD_NAME} #(
    
) (
    input clk, n_rst
);

    

endmodule
